module MAC( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [3:0] io_in_a, // @[:@6.4]
  input  [3:0] io_in_b, // @[:@6.4]
  input  [3:0] io_in_c, // @[:@6.4]
  output [7:0] io_out // @[:@6.4]
);
  wire [7:0] _T_13; // @[combinational_logic.scala 15:22:@8.4]
  wire [7:0] _GEN_0; // @[combinational_logic.scala 15:33:@9.4]
  wire [8:0] _T_14; // @[combinational_logic.scala 15:33:@9.4]
  assign _T_13 = io_in_a * io_in_b; // @[combinational_logic.scala 15:22:@8.4]
  assign _GEN_0 = {{4'd0}, io_in_c}; // @[combinational_logic.scala 15:33:@9.4]
  assign _T_14 = _T_13 + _GEN_0; // @[combinational_logic.scala 15:33:@9.4]
  assign io_out = _T_13 + _GEN_0; // @[combinational_logic.scala 15:10:@11.4]
endmodule
