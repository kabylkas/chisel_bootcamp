module Arbiter( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_fifo_valid, // @[:@6.4]
  output        io_fifo_ready, // @[:@6.4]
  input  [15:0] io_fifo_data, // @[:@6.4]
  output        io_pe0_valid, // @[:@6.4]
  input         io_pe0_ready, // @[:@6.4]
  output [15:0] io_pe0_data, // @[:@6.4]
  output        io_pe1_valid, // @[:@6.4]
  input         io_pe1_ready, // @[:@6.4]
  output [15:0] io_pe1_data // @[:@6.4]
);
  wire  _GEN_3; // @[exercise2.scala 28:25:@13.6]
  assign _GEN_3 = io_pe0_ready ? 1'h0 : io_pe1_ready; // @[exercise2.scala 28:25:@13.6]
  assign io_fifo_ready = io_pe0_ready | io_pe1_ready; // @[exercise2.scala 25:17:@11.4]
  assign io_pe0_valid = io_fifo_valid ? io_pe0_ready : 1'h0; // @[exercise2.scala 29:20:@14.8 exercise2.scala 32:20:@19.10 exercise2.scala 35:20:@23.10 exercise2.scala 39:20:@28.6]
  assign io_pe0_data = io_fifo_data; // @[exercise2.scala 23:15:@8.4]
  assign io_pe1_valid = io_fifo_valid ? _GEN_3 : 1'h0; // @[exercise2.scala 30:20:@15.8 exercise2.scala 33:20:@20.10 exercise2.scala 36:20:@24.10 exercise2.scala 40:20:@29.6]
  assign io_pe1_data = io_fifo_data; // @[exercise2.scala 24:15:@9.4]
endmodule
