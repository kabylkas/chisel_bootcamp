module PolyCircuit( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [1:0]  io_select, // @[:@6.4]
  input  [31:0] io_x, // @[:@6.4]
  output [31:0] io_fofx // @[:@6.4]
);
  wire [63:0] _T_13; // @[exercise1.scala 17:16:@10.4]
  wire [31:0] _GEN_0; // @[exercise1.scala 15:18:@9.4 exercise1.scala 17:8:@11.4]
  wire [31:0] x_sq; // @[exercise1.scala 15:18:@9.4 exercise1.scala 17:8:@11.4]
  wire [35:0] _T_15; // @[exercise1.scala 24:19:@12.4]
  wire [36:0] _T_17; // @[exercise1.scala 24:33:@13.4]
  wire [36:0] _GEN_1; // @[exercise1.scala 24:26:@14.4]
  wire [37:0] _T_18; // @[exercise1.scala 24:26:@14.4]
  wire [36:0] _T_19; // @[exercise1.scala 24:26:@15.4]
  wire [36:0] _T_20; // @[exercise1.scala 24:26:@16.4]
  wire [37:0] _T_22; // @[exercise1.scala 24:40:@17.4]
  wire [36:0] _T_23; // @[exercise1.scala 24:40:@18.4]
  wire [36:0] _T_24; // @[exercise1.scala 24:40:@19.4]
  wire [31:0] _GEN_2; // @[exercise1.scala 14:20:@8.4 exercise1.scala 24:12:@20.4]
  assign _T_13 = $signed(io_x) * $signed(io_x); // @[exercise1.scala 17:16:@10.4]
  assign _GEN_0 = _T_13[31:0]; // @[exercise1.scala 15:18:@9.4 exercise1.scala 17:8:@11.4]
  assign x_sq = $signed(_GEN_0); // @[exercise1.scala 15:18:@9.4 exercise1.scala 17:8:@11.4]
  assign _T_15 = $signed(32'sh4) * $signed(x_sq); // @[exercise1.scala 24:19:@12.4]
  assign _T_17 = $signed(32'sha) * $signed(io_x); // @[exercise1.scala 24:33:@13.4]
  assign _GEN_1 = {{1{_T_15[35]}},_T_15}; // @[exercise1.scala 24:26:@14.4]
  assign _T_18 = $signed(_GEN_1) - $signed(_T_17); // @[exercise1.scala 24:26:@14.4]
  assign _T_19 = $signed(_GEN_1) - $signed(_T_17); // @[exercise1.scala 24:26:@15.4]
  assign _T_20 = $signed(_T_19); // @[exercise1.scala 24:26:@16.4]
  assign _T_22 = $signed(_T_20) - $signed(37'sh5); // @[exercise1.scala 24:40:@17.4]
  assign _T_23 = $signed(_T_20) - $signed(37'sh5); // @[exercise1.scala 24:40:@18.4]
  assign _T_24 = $signed(_T_23); // @[exercise1.scala 24:40:@19.4]
  assign _GEN_2 = _T_24[31:0]; // @[exercise1.scala 14:20:@8.4 exercise1.scala 24:12:@20.4]
  assign io_fofx = $signed(_GEN_2); // @[exercise1.scala 27:11:@21.4]
endmodule
